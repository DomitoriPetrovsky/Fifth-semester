library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


package iir_config is

    constant IIR_ORDER : natural := 7;

    constant IIR_IWL : natural := 16;

    constant IIR_CWL: natural := 20;
    

    type VECTOR_OF_STD_L_V is array (natural range <>) of std_logic_vector(IIR_CWL - 1 downto 0);

    
    
	-----------------------------------------------------------
    --Butter
	-----------------------------------------------------------
    constant COEFFS_A_L : VECTOR_OF_STD_L_V :=
    ( 
    "00001000000000000000",
    "11010110000110110010",
    "01011111011010110000",
    "10000101101110100101",
   "01011111000011111110",
    "11010011001101101001",
    "00001011110101000000",
    "11111110101001100111"
    );

    constant COEFFS_B_L : VECTOR_OF_STD_L_V :=
    (
    "00000000000000000000",
    "00000000000000000001",
    "00000000000000000011",
    "00000000000000000110",
    "00000000000000000110",
    "00000000000000000011",
    "00000000000000000001",
    "00000000000000000000"
    );
	
	-----------------------------------------------------------
	--TEST
	-----------------------------------------------------------
    constant COEFFS_A_T : VECTOR_OF_STD_L_V :=
    ( 
    "00000000000000000000",
    "00000000000000000000",
    "00000000000000000000",
    "00000000000000000000",
    "00000000000000000000",
    "00000000000000000000",
    "00000000000000000000",
    "00000000000000000000"
    );

    constant COEFFS_B_T : VECTOR_OF_STD_L_V :=
    (
    "11111011000000000000",
    "00000001000000000000",
    "11111110000000000000",
    "11111100000000000000",
    "00000100000000000000",
    "00000010000000000000",
    "11111111000000000000",
    "00000101000000000000"
    );
	

	
	constant COEFFS_B : VECTOR_OF_STD_L_V := COEFFS_B_L;
    constant COEFFS_A : VECTOR_OF_STD_L_V := COEFFS_A_T;
end iir_config;

--package body iir_config is
  
--end iir_config;