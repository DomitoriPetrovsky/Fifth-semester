package automat_states is
  
  type fsm_in_type is (z1, z2, z3);
  type fsm_out_type is (w1, w2, w3, o);
end automat_states;
 
package body automat_states is
  
end automat_states;