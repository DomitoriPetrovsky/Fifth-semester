library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


package iir_config is

    constant IIR_ORDER : natural := 7;

    constant IIR_IWL : natural := 16;

    constant IIR_CWL: natural := 20;
    

    type VECTOR_OF_STD_L_V is array (natural range <>) of std_logic_vector(IIR_CWL - 1 downto 0);

    
    
	-----------------------------------------------------------
    --Butter Low
	-----------------------------------------------------------
    constant COEFFS_A_L : VECTOR_OF_STD_L_V :=
    ( 
    "00001000000000000000",
    "11010110000110110010",
    "01011111011010110000",
    "10000101101110100101",
    "01011111000011111110",
    "11010011001101101001",
    "00001011110101000000",
    "11111110101001100111"
    );

    constant COEFFS_B_L : VECTOR_OF_STD_L_V :=
    (
    "00000000000000000000",
    "00000000000000000001",
    "00000000000000000011",
    "00000000000000000110",
    "00000000000000000110",
    "00000000000000000011",
    "00000000000000000001",
    "00000000000000000000"
    );
	
	-----------------------------------------------------------
    --Butter Medium
	-----------------------------------------------------------
	
	--CONSTANT IIR_IWL: NATURAL := 16;
	--CONSTANT IIR_CWL: NATURAL := 28; можно и 26
	
    constant COEFFS_A_M : VECTOR_OF_STD_L_V :=
    ( 
    "0000000000001000000000000000",   
	"1111111110101101000000100110",   
	"0000000110011011110111011100",   
	"1111101011110010011101100111",   
	"0000101100110100011100011011",   
	"1110110101110101011000100111",   
	"0001011110011000110000100010",   
	"1110100010001011110010101011",   
	"0001001001001011001100101000",   
	"1111010011011011000110000010",   
	"0000010100111000101000010010",   
	"1111111000101100101010001001",   
	"0000000001110011011001000110",   
	"1111111111101101111101101000",  
	"0000000000000001010110011001"
    );

    constant COEFFS_B_M : VECTOR_OF_STD_L_V :=
    (
    "0000000000000000000000000000",   
	"0000000000000000000000000000",   
	"1111111111111111111111111111",  
	"0000000000000000000000000000",  
	"0000000000000000000000000011",  
	"0000000000000000000000000000",   
	"1111111111111111111111111010",  
	"0000000000000000000000000000",   
	"0000000000000000000000000110",   
	"0000000000000000000000000000",   
	"1111111111111111111111111101",   
	"0000000000000000000000000000",   
	"0000000000000000000000000001",   
	"0000000000000000000000000000",
	"0000000000000000000000000000"
    );
	
	-----------------------------------------------------------
	--TEST
	-----------------------------------------------------------
    constant COEFFS_A_T_2 : VECTOR_OF_STD_L_V :=
    ( 
    "00000000000000000000",
    "11010110000110110010",
    "01011111011010110000",
    "00000000000000000000",
    "00000000000000000000",
    "00000000000000000000",
    "00000000000000000000",
    "00000000000000000000"
    );

	constant COEFFS_B_T_2 : VECTOR_OF_STD_L_V :=
    (
    "00001000000000000000",
    "00000000000000000000",
    "00000000000000000000",
    "00000000000000000000",
    "00000000000000000000",
    "00000000000000000000",
    "00000000000000000000",
    "00000000000000000000"
    );
	
	constant COEFFS_A_T_1 : VECTOR_OF_STD_L_V :=
    ( 
    "00000000000000000000",
    "00000000000000000000",
    "00000000000000000000",
    "00000000000000000000",
    "00000000000000000000",
    "00000000000000000000",
    "00000000000000000000",
    "00000000000000000000"
    );
	
    constant COEFFS_B_T_1 : VECTOR_OF_STD_L_V :=
    (
    "11111011000000000000",
    "00000001000000000000",
    "11111110000000000000",
    "11111100000000000000",
    "00000100000000000000",
    "00000010000000000000",
    "11111111000000000000",
    "00000101000000000000"
    );
	

	
	constant COEFFS_B : VECTOR_OF_STD_L_V := COEFFS_B_L;
    constant COEFFS_A : VECTOR_OF_STD_L_V := COEFFS_A_L;
end iir_config;

--package body iir_config is
  
--end iir_config;